-- Code your design here
library IEEE;
use IEEE.std_logic_1164.all;

entity mycomponent is
end mycomponent;

architecture myarchitecture of mycomponent is
begin 
end myarchitecture;